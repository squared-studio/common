////////////////////////////////////////////////////////////////////////////////////////////////////
//
//    AUTHOR      : ...
//    EMAIL       : ...
//
//    MODULE      : ...
//    DESCRIPTION : ...
//
////////////////////////////////////////////////////////////////////////////////////////////////////

//`define ENABLE_DUMPFILE

module tb_model;

    ////////////////////////////////////////////////////////////////////////////////////////////////
    // IMPORTS
    ////////////////////////////////////////////////////////////////////////////////////////////////

    // bring in the testbench essentials functions and macros
    `include "tb_essentials.sv"

    ////////////////////////////////////////////////////////////////////////////////////////////////
    // LOCALPARAMS
    ////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////
    // TYPEDEFS
    ////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SIGNALS
    ////////////////////////////////////////////////////////////////////////////////////////////////

    // generates static task start_clk_i with tHigh:3 tLow:7
    `CREATE_CLK(clk_i, 3, 7)

    bit arst_n = 1;

    ////////////////////////////////////////////////////////////////////////////////////////////////
    // VARIABLES
    ////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////
    // INTERFACES
    ////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////
    // CLASSES
    ////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////
    // ASSIGNMENTS
    ////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////
    // RTLS
    ////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////
    // METHODS
    ////////////////////////////////////////////////////////////////////////////////////////////////

    task static apply_reset ();
        #100;
        arst_n = 0;
        #100;
        arst_n = 1;
        #100;
    endtask

    ////////////////////////////////////////////////////////////////////////////////////////////////
    // PROCEDURALS
    ////////////////////////////////////////////////////////////////////////////////////////////////

    initial begin
        apply_reset();
        start_clk_i();

        @ (posedge clk_i);
        result_print (1, "This is a PASS");
        @ (posedge clk_i);
        result_print (0, "And this is a FAIL");

        $finish;

    end

endmodule
