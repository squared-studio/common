// Register file for floating point 
// ### Author : Md. Mohiuddin Reyad (mreyad30207@gmail.com)

module rv_float_reg_file #(
    parameter int FLEN = 32,
    parameter int ELEM_WIDTH = 7
) (
  input  logic                    clk_i,   // Global clock
  input  logic                    arst_ni, // Asynchronous reset
  
  input  logic [$clog2(FLEN)-1:0] rd_addr_i,  // read address 
  input  logic [ELEM_WIDTH -1:0 ] rd_data_i,  //read data
  input  logic                    rd_en_i,   // read enable
  
  input  logic [$clog2(FLEN)-1:0] rs1_addr_i,
  output logic [ELEM_WIDTH -1:0 ] rs1_data_o,
  
  input  logic [$clog2(FLEN)-1:0] rs2_addr_i,
  output logic [ELEM_WIDTH -1:0 ] rs2_data_o,
  
  input  logic [$clog2(FLEN)-1:0] rs3_addr_i,
  output logic [ELEM_WIDTH -1:0 ] rs3_data_o
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENCIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef SIMULATION
  initial begin
    if (DATA_WIDTH > 2) begin
      $display("\033[7;31m%m DATA_WIDTH\033[0m");
    end
  end
`endif  // SIMULATION

endmodule
