// Description here
// ### Author : Walid Akash (walidakash070@gmail.com)

//`include "axi4/typedef.svh"
//`include "axi4/assign.svh"
//`include "axi4l/typedef.svh"
//`include "axi4l/assign.svh"
//`include "vip/bus_dvr_mon.svh"

//`include "vip/string_ops_pkg.sv"

module xbar_tb;

  //`define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  localparam int ElemWidth = 4;
  localparam int NumElem = 6;


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  logic [NumElem-1:0][$clog2(NumElem)-1:0] select_i;
  logic [NumElem-1:0][ElemWidth-1:0] inputs_i;
  logic [NumElem-1:0][ElemWidth-1:0] outputs_o;

  // generates static task start_clk_i with tHigh:3 tLow:7
  //`CREATE_CLK(clk_i, 3, 7)

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  logic error = 0;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  xbar #(
      .ElemWidth(ElemWidth),
      .NumElem  (NumElem)
  ) xbar_dut (
      .select_i (select_i),
      .inputs_i (inputs_i),
      .outputs_o(outputs_o)
  );


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // task static apply_reset();
  //  #5;
  //  arst_ni = 0;
  //  #5;
  //  arst_ni = 1;
  //  #5;
  //endtask

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin
    //apply_reset();
    //start_clk_i();
    for (int i = 0; i < NumElem; i++) begin
      inputs_i[i] = $urandom;
      select_i[i] = $urandom_range(0, NumElem - 1);
    end
    #200;

    $display("inputs_i = %p", inputs_i);
    $display("select_i = %p", select_i);
    $display("outputs_o = %p", outputs_o);

    for (int i = 0; i < NumElem; i++) begin
      if (outputs_o[i] == inputs_i[select_i[i]]) begin
        error++;
      end else begin
        error = error;
      end
    end
    result_print(error == 0, "CrossBar verified");

    $finish;

  end

endmodule
