/*
Description
Author : Foez Ahmed (foez.official@gmail.com)
<br>This file is part of squared-studio:common
<br>Copyright (c) 2024 squared-studio
<br>Licensed under the MIT License
<br>See LICENSE file in the project root for full license information
*/

module shifter_tb;

  //`define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  localparam int DataWidth = 16;
  localparam int ShiftWidth = 3;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns
  `CREATE_CLK(clk_i, 4ns, 6ns)

  logic [ShiftWidth-1:0] shift_i = '0;
  logic                  right_shift_i = '0;
  logic [ DataWidth-1:0] data_i = '0;
  logic [ DataWidth-1:0] data_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  int                    pass = 0;
  int                    fail = 0;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  shifter #(
      .DATA_WIDTH (DataWidth),
      .SHIFT_WIDTH(ShiftWidth)
  ) u_shifter (
      .shift_i(shift_i),
      .right_shift_i(right_shift_i),
      .data_i(data_i),
      .data_o(data_o)
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static rnd_drv();
    fork
      forever begin
        @(posedge clk_i);
        shift_i       <= $urandom;
        right_shift_i <= $urandom;
        data_i        <= $urandom;
      end
    join_none
  endtask

  task static check();
    fork
      forever begin
        logic [DataWidth-1:0] expectation;
        @(posedge clk_i);
        if (right_shift_i) expectation = data_i >> shift_i;
        else expectation = data_i << shift_i;
        if (expectation === data_o) pass++;
        else fail++;
      end
    join_none
  endtask

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    start_clk_i();
    rnd_drv();
    check();

    repeat (50) @(posedge clk_i);
    result_print(!fail, $sformatf("%0d/%0d Passed", pass, pass+fail));

    $finish;

  end

endmodule
