////////////////////////////////////////////////////////////////////////////////////////////////////
//
//    AUTHOR      : ...
//    EMAIL       : ...
//
//    MODULE      : ...
//    DESCRIPTION : ...
//
////////////////////////////////////////////////////////////////////////////////////////////////////

module bin_to_gray_tb;

    ////////////////////////////////////////////////////////////////////////////////////////////////////
    // IMPORTS
    ////////////////////////////////////////////////////////////////////////////////////////////////////

        `include "tb_essentials.sv"

    ////////////////////////////////////////////////////////////////////////////////////////////////////
    // LOCALPARAMS
    ////////////////////////////////////////////////////////////////////////////////////////////////////

        localparam int DataWidth = 4;

    ////////////////////////////////////////////////////////////////////////////////////////////////////
    // TYPEDEFS
    ////////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////////
    // SIGNALS
    ////////////////////////////////////////////////////////////////////////////////////////////////////
        `CREATE_CLK(clk_i, 3, 7)

        bit arst_n = 1;

        logic [DataWidth-1:0] data_in_i;
        logic [DataWidth-1:0] data_out_o;

        logic [DataWidth-1:0] data_out_temp;
        int pass;
        int fail;

    ////////////////////////////////////////////////////////////////////////////////////////////////////
    // INTERFACES
    ////////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////////
    // CLASSES
    ////////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////////
    // ASSIGNMENTS
    ////////////////////////////////////////////////////////////////////////////////////////////////////



    ////////////////////////////////////////////////////////////////////////////////////////////////////
    // RTLS
    ////////////////////////////////////////////////////////////////////////////////////////////////////

        bin_to_gray #(
            .DataWidth (DataWidth)
        ) bin_to_gray_dut (
            .data_in_i  ( data_in_i  ),
            .data_out_o ( data_out_o )
        );

    ////////////////////////////////////////////////////////////////////////////////////////////////////
    // METHODS
    ////////////////////////////////////////////////////////////////////////////////////////////////////
    task static start_clock  ();
        fork
            forever
            begin
                clk_i  = 1; #5;
                clk_i  = 0; #5;
            end
        join_none
    endtask : start_clock

    task static apply_reset ();
        #100;
        arst_n = 0;
        #100;
        arst_n = 1;
        #100;
    endtask

    ////////////////////////////////////////////////////////////////////////////////////////////////////
    // PROCEDURALS
    ////////////////////////////////////////////////////////////////////////////////////////////////////

        initial begin
            $dumpfile("raw.vcd");
            $dumpvars();

            apply_reset();
            start_clock();
            repeat (1) @(posedge clk_i)
            begin
                //data_in_i =$urandom_range(0,15);
                $monitor("Binary = %b  Gray   = %b", data_in_i, data_out_o);
                data_in_i = 4'b0000; #1;
                data_in_i = 4'b0001; #1;
                data_in_i = 4'b0010; #1;
                data_in_i = 4'b0011; #1;
                data_in_i = 4'b0100; #1;
                data_in_i = 4'b0101; #1;
                data_in_i = 4'b0110; #1;
                data_in_i = 4'b0111; #1;
                data_in_i = 4'b1000; #1;
                data_in_i = 4'b1001; #1;
                data_in_i = 4'b1010; #1;
                data_in_i = 4'b1011; #1;
                data_in_i = 4'b1100; #1;
                data_in_i = 4'b1101; #1;
                data_in_i = 4'b1110; #1;
                data_in_i = 4'b1111;

           /*
                for(int i=0;i<15;i++) begin
                assign data_out_temp[i] = data_in_i[i] ^ data_in_i[i+1];
            end
            // $monitor("Binary = %b  Gray   = %b", data_in_i, data_out_o); end
            
            foreach(data_out_o[j]) begin
                if(data_out_temp == data_out_o) begin
                    pass++;
                    result_print (1, "This is a PASS");
                end
                else
                    fail++;
                    result_print (0, "And this is a FAIL");
                    */
            #100;
            $finish;
            end
        end
endmodule
