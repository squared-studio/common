// ### Author : Foez Ahmed (foez.official@gmail.com)

(* no_ungroup *) (* no_boundary_optimization *) (* dont_touch = "true" *)
module buffer #(
    parameter int WIDTH = 8
) (
    input  logic [WIDTH-1:0] d_i,
    output logic [WIDTH-1:0] q_o
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  logic [WIDTH-1:0] mid_wire;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  inverter #(
      .WIDTH(WIDTH)
  ) inverter_in (
      .d_i(d_i),
      .q_o(mid_wire)
  );

  inverter #(
      .WIDTH(WIDTH)
  ) inverter_out (
      .d_i(mid_wire),
      .q_o(q_o)
  );

endmodule
