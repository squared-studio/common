package memory_pkg;

  `include "vip/memory_ops.svh"

  class byte_memory;
    //////////////////////////////////////////////////////////////////////////////////////////////////
    //-SIGNALS
    //////////////////////////////////////////////////////////////////////////////////////////////////

    bit [7:0] mem[longint];

    //////////////////////////////////////////////////////////////////////////////////////////////////
    //-METHODS
    //////////////////////////////////////////////////////////////////////////////////////////////////

    function automatic load_image(input string file);
      `LOAD_HEX(file, mem)
    endfunction

    function automatic save_image(input string file);
      `SAVE_HEX(file, mem)
    endfunction

  endclass

endpackage
