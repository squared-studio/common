// Description here
// ### Author : Foez Ahmed (foez.official@gmail.com)

module uart_if_tb;

  `define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  uart_if u1 ();

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  assign u1.rx = u1.tx;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    u1.set_baud(20000000);
    u1.set_data_width(4);
    u1.set_parity(0);
    u1.set_stop_width(1);

    $display("baud: %0d", u1.get_baud());
    $display("data_width: %0d", u1.get_data_width());
    $display("parity: %0d", u1.get_parity());
    $display("stop_width: %0d", u1.get_stop_width());

    u1.send('hF);
    u1.send('h0);
    u1.send('hE);
    u1.send('h2);

    do #1ns; while (u1.is_tx_active() || u1.is_rx_active());

    $display("GOT:0x%h", u1.recv());
    $display("GOT:0x%h", u1.recv());
    $display("GOT:0x%h", u1.recv());
    $display("GOT:0x%h", u1.recv());

    $finish;

  end

endmodule
