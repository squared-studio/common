// Clock gate
// ### Author : Razu Ahamed(en.razu.ahamed@gmail.com)

module clk_gate (
  input  logic cp ,
  input  logic e  ,
  input  logic te ,
  output logic q
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  logic temp;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  assign q = te?cp:temp;
  and(temp,cp,e);

endmodule
