// A simple encoder module for translating single wires into address and address valid
// ### Author : Foez Ahmed (foez.official@gmail.com)

module encoder #(
    parameter int ADDR_WIDTH = 4  // Code with
) (
    input  logic [2**ADDR_WIDTH-1:0] select_i,     // Wire input
    output logic [   ADDR_WIDTH-1:0] addr_o,       // Address output
    output logic                     addr_valid_o  // Address Valid output
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  wire [ADDR_WIDTH-1:0] addr;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  assign addr_valid_o = |select_i;

  for (genvar i = 0; i < 2 ** ADDR_WIDTH; i++) begin : g_addr
    assign addr = select_i[i] ? i : 'z;
  end

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  for (genvar i = 0; i < ADDR_WIDTH; i++) begin : g_buf_addr_o
    buf (addr_o[i], addr[i]);
  end

endmodule
