// Description
// ### Author : Foez Ahmed (foez.official@gmail.com)

module edge_detector #(
    parameter bit POSEDGE = 1,
    parameter bit NEGEDGE = 1
) (
    input  logic arst_ni,
    input  logic clk_i,
    input  logic d_i,
    output logic posedge_o,
    output logic negedge_o
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  logic q;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  if (POSEDGE) begin : g_pos_assign
    assign posedge_o = d_i & ~q;
  end else begin : g_pos_default
    assign posedge_o = '0;
  end

  if (NEGEDGE) begin : g_neg_assign
    assign negedge_o = ~d_i & q;
  end else begin : g_neg_default
    assign negedge_o = '0;
  end

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENCIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  always_ff @(posedge clk_i or negedge arst_ni) begin
    if (~arst_ni) begin
      q <= '0;
    end else begin
      q <= d_i;
    end
  end

endmodule
