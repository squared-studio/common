// General purpose Encoder
// ### Author : Foez Ahmed (foez.official@gmail.com)

module encoder #(
    parameter int NUM_WIRE = 4  // Number of output wires
) (
    input  logic [        NUM_WIRE-1:0] d_i,          // Wire input
    output logic [$clog2(NUM_WIRE)-1:0] addr_o,       // Address output
    output logic                        addr_valid_o  // Address Valid output
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  wire [$clog2(NUM_WIRE)-1:0] addr;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  assign addr_valid_o = |d_i;

  for (genvar i = 0; i < NUM_WIRE; i++) begin : g_addr
    assign addr = d_i[i] ? i : 'z;
  end

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  for (genvar i = 0; i < $clog2(NUM_WIRE); i++) begin : g_buf_addr_o
    buf (addr_o[i], addr[i]);
  end

endmodule
