package axi4_pkg;

  class axi4_driver #(
    parameter int AddressWidth = 0 
  );
  //`define AXI4_T(__NM__, __AW__, __DW__, __IRW__, __IWW__, __UREQW__, __UDTAW__, __URSPW__)
  endclass

endpackage
