// ### Author : Foez Ahmed (foez.official@gmail.com)

module fixed_priority_arbiter #(
    parameter int NUM_REQ = 4
) (
    input  logic                       allow_req_i,
    input  logic [        NUM_REQ-1:0] req_i,
    output logic [$clog2(NUM_REQ)-1:0] gnt_addr_o,
    output logic                       gnt_addr_valid_o
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  logic addr_valid_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  assign gnt_addr_valid_o = allow_req_i & addr_valid_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  priority_encoder #(
      .NUM_WIRE(NUM_REQ),
      .HIGH_INDEX_PRIORITY(0)
  ) priority_encoder_dut (
      .d_i(req_i),
      .addr_o(gnt_addr_o),
      .addr_valid_o(addr_valid_o)
  );

endmodule
