// Description here
// ### Author : name (email)

//`include "axi4_typedef.svh"
//`include "axi4_assign.svh"
`include "axi4l_typedef.svh"
//`include "axi4l_assign.svh"
//`include "vip/bus_dvr_mon.svh"

//`include "vip/string_ops_pkg.sv"

module axi4l_if_tb;

  `define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  `AXI4L_T(axil, 32, 64)

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns
  `CREATE_CLK(clk_i, 4ns, 6ns)

  bit arst_ni = 1;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  axi4l_if #(
      .req_t (axil_req_t),
      .resp_t(axil_resp_t)
  ) axil_bus_dv (
      .clk_i  (clk_i),
      .arst_ni(arst_ni)
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static apply_reset();
    #100;
    arst_ni = 0;
    #100;
    arst_ni = 1;
    #100;
  endtask

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin

    static int fail;

    fail = 0;
    apply_reset();
    start_clk_i();


    // AW channel transaction test
    repeat (50) begin
      axil_aw_chan_t snd;
      axil_aw_chan_t rcv;
      axil_aw_chan_t mon;
      snd.addr = $urandom;
      snd.prot = $urandom;
      fork
        axil_bus_dv.send_aw(snd);
        axil_bus_dv.recv_aw(rcv);
        axil_bus_dv.look_aw(mon);
      join
      if (snd !== rcv || snd !== mon) fail++;
    end
    result_print(!fail, "AW channel OK");

    // W channel transaction test
    repeat (50) begin
      axil_w_chan_t snd;
      axil_w_chan_t rcv;
      axil_w_chan_t mon;
      snd.data = {$urandom, $urandom};
      snd.strb = $urandom;
      fork
        axil_bus_dv.send_w(snd);
        axil_bus_dv.recv_w(rcv);
        axil_bus_dv.look_w(mon);
      join
      if (snd !== rcv || snd !== mon) fail++;
    end
    result_print(!fail, "W channel OK");

    // B channel transaction test
    repeat (50) begin
      axil_b_chan_t snd;
      axil_b_chan_t rcv;
      axil_b_chan_t mon;
      snd.resp = $urandom;
      fork
        axil_bus_dv.send_b(snd);
        axil_bus_dv.recv_b(rcv);
        axil_bus_dv.look_b(mon);
      join
      if (snd !== rcv || snd !== mon) fail++;
    end
    result_print(!fail, "B channel OK");

    // AR channel transaction test
    repeat (50) begin
      axil_ar_chan_t snd;
      axil_ar_chan_t rcv;
      axil_ar_chan_t mon;
      snd.addr = $urandom;
      snd.prot = $urandom;
      fork
        axil_bus_dv.send_ar(snd);
        axil_bus_dv.recv_ar(rcv);
        axil_bus_dv.look_ar(mon);
      join
      if (snd !== rcv || snd !== mon) fail++;
    end
    result_print(!fail, "AR channel OK");

    // R channel transaction test
    repeat (50) begin
      axil_r_chan_t snd;
      axil_r_chan_t rcv;
      axil_r_chan_t mon;
      snd.data = {$urandom, $urandom};
      snd.resp = $urandom;
      fork
        axil_bus_dv.send_r(snd);
        axil_bus_dv.recv_r(rcv);
        axil_bus_dv.look_r(mon);
      join
      if (snd !== rcv || snd !== mon) fail++;
    end
    result_print(!fail, "R channel OK");

    $finish;

  end

endmodule
