// Clock gate
// ### Author : Foez Ahmed (foez.official@gmail.com)

module clk_gate #(
) (
    input  logic arst_ni,
    input  logic clk_i,
    input  logic en_i,
    output logic clk_o
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  logic dff_out;
  assign clk_o = clk_i & dff_out;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  dual_synchronizer #(
      .FIRST_FF_EDGE_POSEDGED(1),
      .LAST_FF_EDGE_POSEDGED (0)
  ) clk1_ffb2b (
      .clk_i  (clk_i),
      .arst_ni(arst_ni),
      .en_i   ('1),
      .d_i    (en_i),
      .q_o    (dff_out)
  );

endmodule
