module encoder_tb;

  //`define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  localparam int NumWire = 8;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  reg  [        NumWire-1:0] d_i;
  wire [$clog2(NumWire)-1:0] addr_o;
  wire                       addr_valid_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  encoder #(
      .NUM_WIRE(NumWire)
  ) encoder_dut (
      .d_i(d_i),
      .addr_o(addr_o),
      .addr_valid_o(addr_valid_o)
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin

    for (int i = 0; i < 2 ** NumWire; i++) begin
      //d_i = 8'b0100_0000;
      d_i = i;
      #5;
      $display("number of test =%0d, d_i = 0b%b, addr_o = 0b%b addr_valid_o = 0b%b", i, d_i,
               addr_o, addr_valid_o);
    end

    result_print(1, "This is a PASS");

    $finish;

  end
endmodule
